// ============================================================================
//        __
//   \\__/ o\    (C) 2020  Robert Finch, Waterloo
//    \  __ /    All rights reserved.
//     \/_//     robfinch<remove>@finitron.ca
//       ||
//
//	DPD1000Decode.sv
//
// BSD 3-Clause License
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// 1. Redistributions of source code must retain the above copyright notice, this
//    list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright notice,
//    this list of conditions and the following disclaimer in the documentation
//    and/or other materials provided with the distribution.
//
// 3. Neither the name of the copyright holder nor the names of its
//    contributors may be used to endorse or promote products derived from
//    this software without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
// FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
// DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
// OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//                                                                          
// ============================================================================

module DPD1000Decode(clk, i, o);
input clk;
input [9:0] i;
output [11:0] o;

reg [9:0] i1;
genvar g;

(* ram_style="block" *)
reg [11:0] tbl [0:1023];

generate begin : gDPDTbl
for (g = 0; g < 1024; g = g + 1) begin : gdpdtblloop
	initial begin
		tbl[g] = (g % 10) | (((g / 10) & 15) << 4) | (((g/100) & 15) << 8);
	end
end
end
endgenerate

always @(posedge clk)
	i1 <= i;
	
assign o = tbl[i1];

endmodule

module DPDDecodeN(clk, i, o);
parameter N=11;
input clk;
input [N*10-1:0] i;
output [N*12-1:0] o;

genvar g;

generate begin : gDPD
	for (g = 0; g < N; g = g + 1) begin : gdpddloop
		DPD1000Decode(clk, i[g*10+9:g*10], o[g*12+11:g*12]);
	end
end
endgenerate

endmodule
